library ieee;
use ieee.std_logic_1164.all;

entity system_management is
end entity;

architecture arch_system_management of system_management is
begin
end architecture;