library ieee;
use ieee.std_logic_1164.all;

entity add is

end entity;
    port(
        clk : in std_logic;
        input : in std_logic_vector();
        output : out std_logic_vector()
    );
architecture arch_add of add is

begin

end architecture;