library ieee;
use ieee.std_logic_1164.all;

entity registers is

end entity;

architecture arch_registers of registers is

begin

end architecture;