library ieee;
use ieee.std_logic_1164.all;

entity top is
    port(
        clk : in std_logic;
    );
end entity;

architecture arch_top of top is

begin

end architecture;