library ieee;
use ieee.std_logic_1164.all;

entity memory_instruction is

end entity;

architecture arch_memory_instruction of memory_instruction is

begin

end architecture;