library ieee;
use ieee.std_logic_1164.all;

entity mux is

end entity;

architecture arch_mux of mux is

begin

end architecture;