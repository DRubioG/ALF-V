library ieee;
use ieee.std_logic_1164.all;

entity alu is

end entity;

architecture arch_alu of alu is

begin

end architecture;