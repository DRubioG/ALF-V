library ieee;
use ieee.std_logic_1164.all;

entity data_memory is

end entity;

architecture arch_data_memory of data_memory is

begin

end architecture;