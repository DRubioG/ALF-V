library ieee;
use ieee.std_logic_1164.all;

entity PC is

end entity;

architecture arch_PC of PC is

begin

end architecture;