library ieee;
use ieee.std_logic_1164.all;

entity decode is
end entity;

architecture arch_decoder of decode is
begin
end architecture;