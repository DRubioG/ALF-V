library ieee;
use ieee.std_logic_1164.all;

entity fetch is
end entity;

architecture arch_fetch of fetch is
begin
end architecture;