library ieee;
use ieee.std_logic_1164.all;

entity imm_gen is

end entity;

architecture arch_imm_gen of imm_gen is

begin

end architecture;